for tarning 5 
 first give me star so 
 send me message on telegram
 @mehdisavari
my shaba:
IR030180000000005309602139
